module decoder16bit(
		input logic [3:0] IN,
		output logic [15:0] OUT);

	always_comb
		case(IN)
			4'b0000: OUT = 16'b0000000000000001;
			4'b0001: OUT = 16'b0000000000000010;
			4'b0010: OUT = 16'b0000000000000100;
			4'b0011: OUT = 16'b0000000000001000;
			4'b0100: OUT = 16'b0000000000010000;
			4'b0101: OUT = 16'b0000000000100000;
			4'b0110: OUT = 16'b0000000001000000;
			4'b0111: OUT = 16'b0000000010000000;
			4'b1000: OUT = 16'b0000000100000000;
			4'b1001: OUT = 16'b0000001000000000;
			4'b1010: OUT = 16'b0000010000000000;
			4'b1011: OUT = 16'b0000100000000000;
			4'b1100: OUT = 16'b0001000000000000;
			4'b1101: OUT = 16'b0010000000000000;
			4'b1110: OUT = 16'b0100000000000000;
			4'b1111: OUT = 16'b1000000000000000;
			default: OUT = 16'b0000000000000000;
		endcase 

endmodule
